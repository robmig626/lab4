module FSM_mem_w_init(clk, wr_en, mem_addr, wr_data);

endmodule 