module FSM_mem_w_init()

endmodule 